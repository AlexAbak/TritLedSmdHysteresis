* EESchema Netlist Version 1.1 (Spice format) creation date: 27.04.2015 13:45:41

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
U1  Net-_R7-Pad1_ Net-_R1-Pad2_ Net-_R5-Pad1_ Net-_P1-Pad2_ Net-_R3-Pad2_ Net-_R6-Pad1_ Net-_R10-Pad2_ Net-_D1-Pad1_ LM393		
R9  Net-_D1-Pad2_ Net-_R7-Pad1_ 220Ω		
R10  Net-_D2-Pad2_ Net-_R10-Pad2_ 220Ω		
D1  Net-_D1-Pad1_ Net-_D1-Pad2_ -		
D2  Net-_D1-Pad1_ Net-_D2-Pad2_ +		
R3  Net-_D1-Pad1_ Net-_R3-Pad2_ ?Ω		
R4  Net-_R3-Pad2_ Net-_P1-Pad2_ ?Ω		
P1  Net-_D1-Pad1_ Net-_P1-Pad2_ Power		
P2  Net-_P2-Pad1_ In		
R8  Net-_R10-Pad2_ Net-_R3-Pad2_ ?Ω		
R6  Net-_R6-Pad1_ Net-_P2-Pad1_ ?Ω		
R7  Net-_R7-Pad1_ Net-_R5-Pad1_ ?Ω		
R5  Net-_R5-Pad1_ Net-_P2-Pad1_ ?Ω		
R1  Net-_D1-Pad1_ Net-_R1-Pad2_ ?Ω		
R2  Net-_R1-Pad2_ Net-_P1-Pad2_ ?Ω		

.end
